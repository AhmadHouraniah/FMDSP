module dadda
(
  input  [16 : 0] x,
  input  [16 : 0] y,
  output [33 : 0] z0,
  output [33 : 0] z1
);

  wire [16 : 0] P [0 : 16];

  wire [525 : 0] S;
  wire [525 : 0] C;

  assign P[0][0] = (x[0] & y[0]);
  assign P[0][1] = (x[0] & y[1]);
  assign P[0][2] = (x[0] & y[2]);
  assign P[0][3] = (x[0] & y[3]);
  assign P[0][4] = (x[0] & y[4]);
  assign P[0][5] = (x[0] & y[5]);
  assign P[0][6] = (x[0] & y[6]);
  assign P[0][7] = (x[0] & y[7]);
  assign P[0][8] = (x[0] & y[8]);
  assign P[0][9] = (x[0] & y[9]);
  assign P[0][10] = (x[0] & y[10]);
  assign P[0][11] = (x[0] & y[11]);
  assign P[0][12] = (x[0] & y[12]);
  assign P[0][13] = (x[0] & y[13]);
  assign P[0][14] = (x[0] & y[14]);
  assign P[0][15] = (x[0] & y[15]);
  assign P[0][16] = ~(x[0] & y[16]);
  assign P[1][0] = (x[1] & y[0]);
  assign P[1][1] = (x[1] & y[1]);
  assign P[1][2] = (x[1] & y[2]);
  assign P[1][3] = (x[1] & y[3]);
  assign P[1][4] = (x[1] & y[4]);
  assign P[1][5] = (x[1] & y[5]);
  assign P[1][6] = (x[1] & y[6]);
  assign P[1][7] = (x[1] & y[7]);
  assign P[1][8] = (x[1] & y[8]);
  assign P[1][9] = (x[1] & y[9]);
  assign P[1][10] = (x[1] & y[10]);
  assign P[1][11] = (x[1] & y[11]);
  assign P[1][12] = (x[1] & y[12]);
  assign P[1][13] = (x[1] & y[13]);
  assign P[1][14] = (x[1] & y[14]);
  assign P[1][15] = (x[1] & y[15]);
  assign P[1][16] = ~(x[1] & y[16]);
  assign P[2][0] = (x[2] & y[0]);
  assign P[2][1] = (x[2] & y[1]);
  assign P[2][2] = (x[2] & y[2]);
  assign P[2][3] = (x[2] & y[3]);
  assign P[2][4] = (x[2] & y[4]);
  assign P[2][5] = (x[2] & y[5]);
  assign P[2][6] = (x[2] & y[6]);
  assign P[2][7] = (x[2] & y[7]);
  assign P[2][8] = (x[2] & y[8]);
  assign P[2][9] = (x[2] & y[9]);
  assign P[2][10] = (x[2] & y[10]);
  assign P[2][11] = (x[2] & y[11]);
  assign P[2][12] = (x[2] & y[12]);
  assign P[2][13] = (x[2] & y[13]);
  assign P[2][14] = (x[2] & y[14]);
  assign P[2][15] = (x[2] & y[15]);
  assign P[2][16] = ~(x[2] & y[16]);
  assign P[3][0] = (x[3] & y[0]);
  assign P[3][1] = (x[3] & y[1]);
  assign P[3][2] = (x[3] & y[2]);
  assign P[3][3] = (x[3] & y[3]);
  assign P[3][4] = (x[3] & y[4]);
  assign P[3][5] = (x[3] & y[5]);
  assign P[3][6] = (x[3] & y[6]);
  assign P[3][7] = (x[3] & y[7]);
  assign P[3][8] = (x[3] & y[8]);
  assign P[3][9] = (x[3] & y[9]);
  assign P[3][10] = (x[3] & y[10]);
  assign P[3][11] = (x[3] & y[11]);
  assign P[3][12] = (x[3] & y[12]);
  assign P[3][13] = (x[3] & y[13]);
  assign P[3][14] = (x[3] & y[14]);
  assign P[3][15] = (x[3] & y[15]);
  assign P[3][16] = ~(x[3] & y[16]);
  assign P[4][0] = (x[4] & y[0]);
  assign P[4][1] = (x[4] & y[1]);
  assign P[4][2] = (x[4] & y[2]);
  assign P[4][3] = (x[4] & y[3]);
  assign P[4][4] = (x[4] & y[4]);
  assign P[4][5] = (x[4] & y[5]);
  assign P[4][6] = (x[4] & y[6]);
  assign P[4][7] = (x[4] & y[7]);
  assign P[4][8] = (x[4] & y[8]);
  assign P[4][9] = (x[4] & y[9]);
  assign P[4][10] = (x[4] & y[10]);
  assign P[4][11] = (x[4] & y[11]);
  assign P[4][12] = (x[4] & y[12]);
  assign P[4][13] = (x[4] & y[13]);
  assign P[4][14] = (x[4] & y[14]);
  assign P[4][15] = (x[4] & y[15]);
  assign P[4][16] = ~(x[4] & y[16]);
  assign P[5][0] = (x[5] & y[0]);
  assign P[5][1] = (x[5] & y[1]);
  assign P[5][2] = (x[5] & y[2]);
  assign P[5][3] = (x[5] & y[3]);
  assign P[5][4] = (x[5] & y[4]);
  assign P[5][5] = (x[5] & y[5]);
  assign P[5][6] = (x[5] & y[6]);
  assign P[5][7] = (x[5] & y[7]);
  assign P[5][8] = (x[5] & y[8]);
  assign P[5][9] = (x[5] & y[9]);
  assign P[5][10] = (x[5] & y[10]);
  assign P[5][11] = (x[5] & y[11]);
  assign P[5][12] = (x[5] & y[12]);
  assign P[5][13] = (x[5] & y[13]);
  assign P[5][14] = (x[5] & y[14]);
  assign P[5][15] = (x[5] & y[15]);
  assign P[5][16] = ~(x[5] & y[16]);
  assign P[6][0] = (x[6] & y[0]);
  assign P[6][1] = (x[6] & y[1]);
  assign P[6][2] = (x[6] & y[2]);
  assign P[6][3] = (x[6] & y[3]);
  assign P[6][4] = (x[6] & y[4]);
  assign P[6][5] = (x[6] & y[5]);
  assign P[6][6] = (x[6] & y[6]);
  assign P[6][7] = (x[6] & y[7]);
  assign P[6][8] = (x[6] & y[8]);
  assign P[6][9] = (x[6] & y[9]);
  assign P[6][10] = (x[6] & y[10]);
  assign P[6][11] = (x[6] & y[11]);
  assign P[6][12] = (x[6] & y[12]);
  assign P[6][13] = (x[6] & y[13]);
  assign P[6][14] = (x[6] & y[14]);
  assign P[6][15] = (x[6] & y[15]);
  assign P[6][16] = ~(x[6] & y[16]);
  assign P[7][0] = (x[7] & y[0]);
  assign P[7][1] = (x[7] & y[1]);
  assign P[7][2] = (x[7] & y[2]);
  assign P[7][3] = (x[7] & y[3]);
  assign P[7][4] = (x[7] & y[4]);
  assign P[7][5] = (x[7] & y[5]);
  assign P[7][6] = (x[7] & y[6]);
  assign P[7][7] = (x[7] & y[7]);
  assign P[7][8] = (x[7] & y[8]);
  assign P[7][9] = (x[7] & y[9]);
  assign P[7][10] = (x[7] & y[10]);
  assign P[7][11] = (x[7] & y[11]);
  assign P[7][12] = (x[7] & y[12]);
  assign P[7][13] = (x[7] & y[13]);
  assign P[7][14] = (x[7] & y[14]);
  assign P[7][15] = (x[7] & y[15]);
  assign P[7][16] = ~(x[7] & y[16]);
  assign P[8][0] = (x[8] & y[0]);
  assign P[8][1] = (x[8] & y[1]);
  assign P[8][2] = (x[8] & y[2]);
  assign P[8][3] = (x[8] & y[3]);
  assign P[8][4] = (x[8] & y[4]);
  assign P[8][5] = (x[8] & y[5]);
  assign P[8][6] = (x[8] & y[6]);
  assign P[8][7] = (x[8] & y[7]);
  assign P[8][8] = (x[8] & y[8]);
  assign P[8][9] = (x[8] & y[9]);
  assign P[8][10] = (x[8] & y[10]);
  assign P[8][11] = (x[8] & y[11]);
  assign P[8][12] = (x[8] & y[12]);
  assign P[8][13] = (x[8] & y[13]);
  assign P[8][14] = (x[8] & y[14]);
  assign P[8][15] = (x[8] & y[15]);
  assign P[8][16] = ~(x[8] & y[16]);
  assign P[9][0] = (x[9] & y[0]);
  assign P[9][1] = (x[9] & y[1]);
  assign P[9][2] = (x[9] & y[2]);
  assign P[9][3] = (x[9] & y[3]);
  assign P[9][4] = (x[9] & y[4]);
  assign P[9][5] = (x[9] & y[5]);
  assign P[9][6] = (x[9] & y[6]);
  assign P[9][7] = (x[9] & y[7]);
  assign P[9][8] = (x[9] & y[8]);
  assign P[9][9] = (x[9] & y[9]);
  assign P[9][10] = (x[9] & y[10]);
  assign P[9][11] = (x[9] & y[11]);
  assign P[9][12] = (x[9] & y[12]);
  assign P[9][13] = (x[9] & y[13]);
  assign P[9][14] = (x[9] & y[14]);
  assign P[9][15] = (x[9] & y[15]);
  assign P[9][16] = ~(x[9] & y[16]);
  assign P[10][0] = (x[10] & y[0]);
  assign P[10][1] = (x[10] & y[1]);
  assign P[10][2] = (x[10] & y[2]);
  assign P[10][3] = (x[10] & y[3]);
  assign P[10][4] = (x[10] & y[4]);
  assign P[10][5] = (x[10] & y[5]);
  assign P[10][6] = (x[10] & y[6]);
  assign P[10][7] = (x[10] & y[7]);
  assign P[10][8] = (x[10] & y[8]);
  assign P[10][9] = (x[10] & y[9]);
  assign P[10][10] = (x[10] & y[10]);
  assign P[10][11] = (x[10] & y[11]);
  assign P[10][12] = (x[10] & y[12]);
  assign P[10][13] = (x[10] & y[13]);
  assign P[10][14] = (x[10] & y[14]);
  assign P[10][15] = (x[10] & y[15]);
  assign P[10][16] = ~(x[10] & y[16]);
  assign P[11][0] = (x[11] & y[0]);
  assign P[11][1] = (x[11] & y[1]);
  assign P[11][2] = (x[11] & y[2]);
  assign P[11][3] = (x[11] & y[3]);
  assign P[11][4] = (x[11] & y[4]);
  assign P[11][5] = (x[11] & y[5]);
  assign P[11][6] = (x[11] & y[6]);
  assign P[11][7] = (x[11] & y[7]);
  assign P[11][8] = (x[11] & y[8]);
  assign P[11][9] = (x[11] & y[9]);
  assign P[11][10] = (x[11] & y[10]);
  assign P[11][11] = (x[11] & y[11]);
  assign P[11][12] = (x[11] & y[12]);
  assign P[11][13] = (x[11] & y[13]);
  assign P[11][14] = (x[11] & y[14]);
  assign P[11][15] = (x[11] & y[15]);
  assign P[11][16] = ~(x[11] & y[16]);
  assign P[12][0] = (x[12] & y[0]);
  assign P[12][1] = (x[12] & y[1]);
  assign P[12][2] = (x[12] & y[2]);
  assign P[12][3] = (x[12] & y[3]);
  assign P[12][4] = (x[12] & y[4]);
  assign P[12][5] = (x[12] & y[5]);
  assign P[12][6] = (x[12] & y[6]);
  assign P[12][7] = (x[12] & y[7]);
  assign P[12][8] = (x[12] & y[8]);
  assign P[12][9] = (x[12] & y[9]);
  assign P[12][10] = (x[12] & y[10]);
  assign P[12][11] = (x[12] & y[11]);
  assign P[12][12] = (x[12] & y[12]);
  assign P[12][13] = (x[12] & y[13]);
  assign P[12][14] = (x[12] & y[14]);
  assign P[12][15] = (x[12] & y[15]);
  assign P[12][16] = ~(x[12] & y[16]);
  assign P[13][0] = (x[13] & y[0]);
  assign P[13][1] = (x[13] & y[1]);
  assign P[13][2] = (x[13] & y[2]);
  assign P[13][3] = (x[13] & y[3]);
  assign P[13][4] = (x[13] & y[4]);
  assign P[13][5] = (x[13] & y[5]);
  assign P[13][6] = (x[13] & y[6]);
  assign P[13][7] = (x[13] & y[7]);
  assign P[13][8] = (x[13] & y[8]);
  assign P[13][9] = (x[13] & y[9]);
  assign P[13][10] = (x[13] & y[10]);
  assign P[13][11] = (x[13] & y[11]);
  assign P[13][12] = (x[13] & y[12]);
  assign P[13][13] = (x[13] & y[13]);
  assign P[13][14] = (x[13] & y[14]);
  assign P[13][15] = (x[13] & y[15]);
  assign P[13][16] = ~(x[13] & y[16]);
  assign P[14][0] = (x[14] & y[0]);
  assign P[14][1] = (x[14] & y[1]);
  assign P[14][2] = (x[14] & y[2]);
  assign P[14][3] = (x[14] & y[3]);
  assign P[14][4] = (x[14] & y[4]);
  assign P[14][5] = (x[14] & y[5]);
  assign P[14][6] = (x[14] & y[6]);
  assign P[14][7] = (x[14] & y[7]);
  assign P[14][8] = (x[14] & y[8]);
  assign P[14][9] = (x[14] & y[9]);
  assign P[14][10] = (x[14] & y[10]);
  assign P[14][11] = (x[14] & y[11]);
  assign P[14][12] = (x[14] & y[12]);
  assign P[14][13] = (x[14] & y[13]);
  assign P[14][14] = (x[14] & y[14]);
  assign P[14][15] = (x[14] & y[15]);
  assign P[14][16] = ~(x[14] & y[16]);
  assign P[15][0] = (x[15] & y[0]);
  assign P[15][1] = (x[15] & y[1]);
  assign P[15][2] = (x[15] & y[2]);
  assign P[15][3] = (x[15] & y[3]);
  assign P[15][4] = (x[15] & y[4]);
  assign P[15][5] = (x[15] & y[5]);
  assign P[15][6] = (x[15] & y[6]);
  assign P[15][7] = (x[15] & y[7]);
  assign P[15][8] = (x[15] & y[8]);
  assign P[15][9] = (x[15] & y[9]);
  assign P[15][10] = (x[15] & y[10]);
  assign P[15][11] = (x[15] & y[11]);
  assign P[15][12] = (x[15] & y[12]);
  assign P[15][13] = (x[15] & y[13]);
  assign P[15][14] = (x[15] & y[14]);
  assign P[15][15] = (x[15] & y[15]);
  assign P[15][16] = ~(x[15] & y[16]);
  assign P[16][0] = ~(x[16] & y[0]);
  assign P[16][1] = ~(x[16] & y[1]);
  assign P[16][2] = ~(x[16] & y[2]);
  assign P[16][3] = ~(x[16] & y[3]);
  assign P[16][4] = ~(x[16] & y[4]);
  assign P[16][5] = ~(x[16] & y[5]);
  assign P[16][6] = ~(x[16] & y[6]);
  assign P[16][7] = ~(x[16] & y[7]);
  assign P[16][8] = ~(x[16] & y[8]);
  assign P[16][9] = ~(x[16] & y[9]);
  assign P[16][10] = ~(x[16] & y[10]);
  assign P[16][11] = ~(x[16] & y[11]);
  assign P[16][12] = ~(x[16] & y[12]);
  assign P[16][13] = ~(x[16] & y[13]);
  assign P[16][14] = ~(x[16] & y[14]);
  assign P[16][15] = ~(x[16] & y[15]);
  assign P[16][16] = (x[16] & y[16]);

  ha HA_00000000 (P[1][16],P[2][15],S[0],C[0]);
  fa FA_00000001 (P[0][16],P[1][15],P[2][14],S[1],C[1]);
  fa FA_00000002 (P[0][15],P[1][14],P[2][13],S[2],C[2]);
  fa FA_00000003 (P[0][14],P[1][13],P[2][12],S[3],C[3]);
  fa FA_00000004 (P[0][13],P[1][12],P[2][11],S[4],C[4]);
  fa FA_00000005 (P[0][12],P[1][11],P[2][10],S[5],C[5]);
  fa FA_00000006 (P[0][11],P[1][10],P[2][9],S[6],C[6]);
  fa FA_00000007 (P[0][10],P[1][9],P[2][8],S[7],C[7]);
  fa FA_00000008 (P[0][9],P[1][8],P[2][7],S[8],C[8]);
  fa FA_00000009 (P[0][8],P[1][7],P[2][6],S[9],C[9]);
  fa FA_00000010 (P[0][7],P[1][6],P[2][5],S[10],C[10]);
  fa FA_00000011 (P[0][6],P[1][5],P[2][4],S[11],C[11]);
  fa FA_00000012 (P[0][5],P[1][4],P[2][3],S[12],C[12]);
  fa FA_00000013 (P[0][4],P[1][3],P[2][2],S[13],C[13]);
  fa FA_00000014 (P[0][3],P[1][2],P[2][1],S[14],C[14]);
  fa FA_00000015 (P[0][2],P[1][1],P[2][0],S[15],C[15]);
  ha HA_00000016 (P[0][1],P[1][0],S[16],C[16]);
  ha HA_00000017 (P[4][16],P[5][15],S[17],C[17]);
  fa FA_00000018 (P[3][16],P[4][15],P[5][14],S[18],C[18]);
  fa FA_00000019 (P[3][15],P[4][14],P[5][13],S[19],C[19]);
  fa FA_00000020 (P[3][14],P[4][13],P[5][12],S[20],C[20]);
  fa FA_00000021 (P[3][13],P[4][12],P[5][11],S[21],C[21]);
  fa FA_00000022 (P[3][12],P[4][11],P[5][10],S[22],C[22]);
  fa FA_00000023 (P[3][11],P[4][10],P[5][9],S[23],C[23]);
  fa FA_00000024 (P[3][10],P[4][9],P[5][8],S[24],C[24]);
  fa FA_00000025 (P[3][9],P[4][8],P[5][7],S[25],C[25]);
  fa FA_00000026 (P[3][8],P[4][7],P[5][6],S[26],C[26]);
  fa FA_00000027 (P[3][7],P[4][6],P[5][5],S[27],C[27]);
  fa FA_00000028 (P[3][6],P[4][5],P[5][4],S[28],C[28]);
  fa FA_00000029 (P[3][5],P[4][4],P[5][3],S[29],C[29]);
  fa FA_00000030 (P[3][4],P[4][3],P[5][2],S[30],C[30]);
  fa FA_00000031 (P[3][3],P[4][2],P[5][1],S[31],C[31]);
  fa FA_00000032 (P[3][2],P[4][1],P[5][0],S[32],C[32]);
  ha HA_00000033 (P[3][1],P[4][0],S[33],C[33]);
  ha HA_00000034 (P[7][16],P[8][15],S[34],C[34]);
  fa FA_00000035 (P[6][16],P[7][15],P[8][14],S[35],C[35]);
  fa FA_00000036 (P[6][15],P[7][14],P[8][13],S[36],C[36]);
  fa FA_00000037 (P[6][14],P[7][13],P[8][12],S[37],C[37]);
  fa FA_00000038 (P[6][13],P[7][12],P[8][11],S[38],C[38]);
  fa FA_00000039 (P[6][12],P[7][11],P[8][10],S[39],C[39]);
  fa FA_00000040 (P[6][11],P[7][10],P[8][9],S[40],C[40]);
  fa FA_00000041 (P[6][10],P[7][9],P[8][8],S[41],C[41]);
  fa FA_00000042 (P[6][9],P[7][8],P[8][7],S[42],C[42]);
  fa FA_00000043 (P[6][8],P[7][7],P[8][6],S[43],C[43]);
  fa FA_00000044 (P[6][7],P[7][6],P[8][5],S[44],C[44]);
  fa FA_00000045 (P[6][6],P[7][5],P[8][4],S[45],C[45]);
  fa FA_00000046 (P[6][5],P[7][4],P[8][3],S[46],C[46]);
  fa FA_00000047 (P[6][4],P[7][3],P[8][2],S[47],C[47]);
  fa FA_00000048 (P[6][3],P[7][2],P[8][1],S[48],C[48]);
  fa FA_00000049 (P[6][2],P[7][1],P[8][0],S[49],C[49]);
  ha HA_00000050 (P[6][1],P[7][0],S[50],C[50]);
  ha HA_00000051 (P[10][16],P[11][15],S[51],C[51]);
  fa FA_00000052 (P[9][16],P[10][15],P[11][14],S[52],C[52]);
  fa FA_00000053 (P[9][15],P[10][14],P[11][13],S[53],C[53]);
  fa FA_00000054 (P[9][14],P[10][13],P[11][12],S[54],C[54]);
  fa FA_00000055 (P[9][13],P[10][12],P[11][11],S[55],C[55]);
  fa FA_00000056 (P[9][12],P[10][11],P[11][10],S[56],C[56]);
  fa FA_00000057 (P[9][11],P[10][10],P[11][9],S[57],C[57]);
  fa FA_00000058 (P[9][10],P[10][9],P[11][8],S[58],C[58]);
  fa FA_00000059 (P[9][9],P[10][8],P[11][7],S[59],C[59]);
  fa FA_00000060 (P[9][8],P[10][7],P[11][6],S[60],C[60]);
  fa FA_00000061 (P[9][7],P[10][6],P[11][5],S[61],C[61]);
  fa FA_00000062 (P[9][6],P[10][5],P[11][4],S[62],C[62]);
  fa FA_00000063 (P[9][5],P[10][4],P[11][3],S[63],C[63]);
  fa FA_00000064 (P[9][4],P[10][3],P[11][2],S[64],C[64]);
  fa FA_00000065 (P[9][3],P[10][2],P[11][1],S[65],C[65]);
  fa FA_00000066 (P[9][2],P[10][1],P[11][0],S[66],C[66]);
  ha HA_00000067 (P[9][1],P[10][0],S[67],C[67]);
  ha HA_00000068 (P[13][16],P[14][15],S[68],C[68]);
  fa FA_00000069 (P[12][16],P[13][15],P[14][14],S[69],C[69]);
  fa FA_00000070 (P[12][15],P[13][14],P[14][13],S[70],C[70]);
  fa FA_00000071 (P[12][14],P[13][13],P[14][12],S[71],C[71]);
  fa FA_00000072 (P[12][13],P[13][12],P[14][11],S[72],C[72]);
  fa FA_00000073 (P[12][12],P[13][11],P[14][10],S[73],C[73]);
  fa FA_00000074 (P[12][11],P[13][10],P[14][9],S[74],C[74]);
  fa FA_00000075 (P[12][10],P[13][9],P[14][8],S[75],C[75]);
  fa FA_00000076 (P[12][9],P[13][8],P[14][7],S[76],C[76]);
  fa FA_00000077 (P[12][8],P[13][7],P[14][6],S[77],C[77]);
  fa FA_00000078 (P[12][7],P[13][6],P[14][5],S[78],C[78]);
  fa FA_00000079 (P[12][6],P[13][5],P[14][4],S[79],C[79]);
  fa FA_00000080 (P[12][5],P[13][4],P[14][3],S[80],C[80]);
  fa FA_00000081 (P[12][4],P[13][3],P[14][2],S[81],C[81]);
  fa FA_00000082 (P[12][3],P[13][2],P[14][1],S[82],C[82]);
  fa FA_00000083 (P[12][2],P[13][1],P[14][0],S[83],C[83]);
  ha HA_00000084 (P[12][1],P[13][0],S[84],C[84]);
  fa FA_00000085 (P[2][16],C[0],S[19],S[85],C[85]);
  fa FA_00000086 (S[0],C[1],S[20],S[86],C[86]);
  fa FA_00000087 (S[1],C[2],S[21],S[87],C[87]);
  fa FA_00000088 (S[2],C[3],S[22],S[88],C[88]);
  fa FA_00000089 (S[3],C[4],S[23],S[89],C[89]);
  fa FA_00000090 (S[4],C[5],S[24],S[90],C[90]);
  fa FA_00000091 (S[5],C[6],S[25],S[91],C[91]);
  fa FA_00000092 (S[6],C[7],S[26],S[92],C[92]);
  fa FA_00000093 (S[7],C[8],S[27],S[93],C[93]);
  fa FA_00000094 (S[8],C[9],S[28],S[94],C[94]);
  fa FA_00000095 (S[9],C[10],S[29],S[95],C[95]);
  fa FA_00000096 (S[10],C[11],S[30],S[96],C[96]);
  fa FA_00000097 (S[11],C[12],S[31],S[97],C[97]);
  fa FA_00000098 (S[12],C[13],S[32],S[98],C[98]);
  fa FA_00000099 (S[13],C[14],S[33],S[99],C[99]);
  fa FA_00000100 (S[14],C[15],P[3][0],S[100],C[100]);
  ha HA_00000101 (S[15],C[16],S[101],C[101]);
  ha HA_00000102 (P[8][16],C[34],S[102],C[102]);
  ha HA_00000103 (S[34],C[35],S[103],C[103]);
  ha HA_00000104 (S[35],C[36],S[104],C[104]);
  fa FA_00000105 (C[17],S[36],C[37],S[105],C[105]);
  fa FA_00000106 (C[18],S[37],C[38],S[106],C[106]);
  fa FA_00000107 (C[19],S[38],C[39],S[107],C[107]);
  fa FA_00000108 (C[20],S[39],C[40],S[108],C[108]);
  fa FA_00000109 (C[21],S[40],C[41],S[109],C[109]);
  fa FA_00000110 (C[22],S[41],C[42],S[110],C[110]);
  fa FA_00000111 (C[23],S[42],C[43],S[111],C[111]);
  fa FA_00000112 (C[24],S[43],C[44],S[112],C[112]);
  fa FA_00000113 (C[25],S[44],C[45],S[113],C[113]);
  fa FA_00000114 (C[26],S[45],C[46],S[114],C[114]);
  fa FA_00000115 (C[27],S[46],C[47],S[115],C[115]);
  fa FA_00000116 (C[28],S[47],C[48],S[116],C[116]);
  fa FA_00000117 (C[29],S[48],C[49],S[117],C[117]);
  fa FA_00000118 (C[30],S[49],C[50],S[118],C[118]);
  ha HA_00000119 (C[31],S[50],S[119],C[119]);
  ha HA_00000120 (C[32],P[6][0],S[120],C[120]);
  fa FA_00000121 (P[11][16],C[51],S[70],S[121],C[121]);
  fa FA_00000122 (S[51],C[52],S[71],S[122],C[122]);
  fa FA_00000123 (S[52],C[53],S[72],S[123],C[123]);
  fa FA_00000124 (S[53],C[54],S[73],S[124],C[124]);
  fa FA_00000125 (S[54],C[55],S[74],S[125],C[125]);
  fa FA_00000126 (S[55],C[56],S[75],S[126],C[126]);
  fa FA_00000127 (S[56],C[57],S[76],S[127],C[127]);
  fa FA_00000128 (S[57],C[58],S[77],S[128],C[128]);
  fa FA_00000129 (S[58],C[59],S[78],S[129],C[129]);
  fa FA_00000130 (S[59],C[60],S[79],S[130],C[130]);
  fa FA_00000131 (S[60],C[61],S[80],S[131],C[131]);
  fa FA_00000132 (S[61],C[62],S[81],S[132],C[132]);
  fa FA_00000133 (S[62],C[63],S[82],S[133],C[133]);
  fa FA_00000134 (S[63],C[64],S[83],S[134],C[134]);
  fa FA_00000135 (S[64],C[65],S[84],S[135],C[135]);
  fa FA_00000136 (S[65],C[66],P[12][0],S[136],C[136]);
  ha HA_00000137 (S[66],C[67],S[137],C[137]);
  ha HA_00000138 (P[15][16],P[16][15],S[138],C[138]);
  fa FA_00000139 (C[68],P[15][15],P[16][14],S[139],C[139]);
  fa FA_00000140 (C[69],P[15][14],P[16][13],S[140],C[140]);
  fa FA_00000141 (C[70],P[15][13],P[16][12],S[141],C[141]);
  fa FA_00000142 (C[71],P[15][12],P[16][11],S[142],C[142]);
  fa FA_00000143 (C[72],P[15][11],P[16][10],S[143],C[143]);
  fa FA_00000144 (C[73],P[15][10],P[16][9],S[144],C[144]);
  fa FA_00000145 (C[74],P[15][9],P[16][8],S[145],C[145]);
  fa FA_00000146 (C[75],P[15][8],P[16][7],S[146],C[146]);
  fa FA_00000147 (C[76],P[15][7],P[16][6],S[147],C[147]);
  fa FA_00000148 (C[77],P[15][6],P[16][5],S[148],C[148]);
  fa FA_00000149 (C[78],P[15][5],P[16][4],S[149],C[149]);
  fa FA_00000150 (C[79],P[15][4],P[16][3],S[150],C[150]);
  fa FA_00000151 (C[80],P[15][3],P[16][2],S[151],C[151]);
  fa FA_00000152 (C[81],P[15][2],P[16][1],S[152],C[152]);
  fa FA_00000153 (C[82],P[15][1],P[16][0],S[153],C[153]);
  ha HA_00000154 (C[83],P[15][0],S[154],C[154]);
  ha HA_00000155 (P[5][16],S[105],S[155],C[155]);
  ha HA_00000156 (S[17],S[106],S[156],C[156]);
  fa FA_00000157 (S[18],C[85],S[107],S[157],C[157]);
  fa FA_00000158 (S[85],C[86],S[108],S[158],C[158]);
  fa FA_00000159 (S[86],C[87],S[109],S[159],C[159]);
  fa FA_00000160 (S[87],C[88],S[110],S[160],C[160]);
  fa FA_00000161 (S[88],C[89],S[111],S[161],C[161]);
  fa FA_00000162 (S[89],C[90],S[112],S[162],C[162]);
  fa FA_00000163 (S[90],C[91],S[113],S[163],C[163]);
  fa FA_00000164 (S[91],C[92],S[114],S[164],C[164]);
  fa FA_00000165 (S[92],C[93],S[115],S[165],C[165]);
  fa FA_00000166 (S[93],C[94],S[116],S[166],C[166]);
  fa FA_00000167 (S[94],C[95],S[117],S[167],C[167]);
  fa FA_00000168 (S[95],C[96],S[118],S[168],C[168]);
  fa FA_00000169 (S[96],C[97],S[119],S[169],C[169]);
  fa FA_00000170 (S[97],C[98],S[120],S[170],C[170]);
  fa FA_00000171 (S[98],C[99],C[33],S[171],C[171]);
  ha HA_00000172 (S[99],C[100],S[172],C[172]);
  ha HA_00000173 (S[100],C[101],S[173],C[173]);
  ha HA_00000174 (S[69],C[121],S[174],C[174]);
  ha HA_00000175 (S[121],C[122],S[175],C[175]);
  ha HA_00000176 (S[122],C[123],S[176],C[176]);
  fa FA_00000177 (C[102],S[123],C[124],S[177],C[177]);
  fa FA_00000178 (C[103],S[124],C[125],S[178],C[178]);
  fa FA_00000179 (C[104],S[125],C[126],S[179],C[179]);
  fa FA_00000180 (C[105],S[126],C[127],S[180],C[180]);
  fa FA_00000181 (C[106],S[127],C[128],S[181],C[181]);
  fa FA_00000182 (C[107],S[128],C[129],S[182],C[182]);
  fa FA_00000183 (C[108],S[129],C[130],S[183],C[183]);
  fa FA_00000184 (C[109],S[130],C[131],S[184],C[184]);
  fa FA_00000185 (C[110],S[131],C[132],S[185],C[185]);
  fa FA_00000186 (C[111],S[132],C[133],S[186],C[186]);
  fa FA_00000187 (C[112],S[133],C[134],S[187],C[187]);
  fa FA_00000188 (C[113],S[134],C[135],S[188],C[188]);
  fa FA_00000189 (C[114],S[135],C[136],S[189],C[189]);
  fa FA_00000190 (C[115],S[136],C[137],S[190],C[190]);
  ha HA_00000191 (C[116],S[137],S[191],C[191]);
  ha HA_00000192 (C[117],S[67],S[192],C[192]);
  ha HA_00000193 (C[118],P[9][0],S[193],C[193]);
  ha HA_00000194 (S[102],S[178],S[194],C[194]);
  ha HA_00000195 (S[103],S[179],S[195],C[195]);
  fa FA_00000196 (S[104],C[155],S[180],S[196],C[196]);
  fa FA_00000197 (S[155],C[156],S[181],S[197],C[197]);
  fa FA_00000198 (S[156],C[157],S[182],S[198],C[198]);
  fa FA_00000199 (S[157],C[158],S[183],S[199],C[199]);
  fa FA_00000200 (S[158],C[159],S[184],S[200],C[200]);
  fa FA_00000201 (S[159],C[160],S[185],S[201],C[201]);
  fa FA_00000202 (S[160],C[161],S[186],S[202],C[202]);
  fa FA_00000203 (S[161],C[162],S[187],S[203],C[203]);
  fa FA_00000204 (S[162],C[163],S[188],S[204],C[204]);
  fa FA_00000205 (S[163],C[164],S[189],S[205],C[205]);
  fa FA_00000206 (S[164],C[165],S[190],S[206],C[206]);
  fa FA_00000207 (S[165],C[166],S[191],S[207],C[207]);
  fa FA_00000208 (S[166],C[167],S[192],S[208],C[208]);
  fa FA_00000209 (S[167],C[168],S[193],S[209],C[209]);
  fa FA_00000210 (S[168],C[169],C[119],S[210],C[210]);
  fa FA_00000211 (S[169],C[170],C[120],S[211],C[211]);
  ha HA_00000212 (S[170],C[171],S[212],C[212]);
  ha HA_00000213 (S[171],C[172],S[213],C[213]);
  ha HA_00000214 (S[172],C[173],S[214],C[214]);
  ha HA_00000215 (P[16][16],C[138],S[215],C[215]);
  ha HA_00000216 (S[138],C[139],S[216],C[216]);
  fa FA_00000217 (P[14][16],S[139],C[140],S[217],C[217]);
  fa FA_00000218 (C[174],S[140],C[141],S[218],C[218]);
  fa FA_00000219 (C[175],S[141],C[142],S[219],C[219]);
  fa FA_00000220 (C[176],S[142],C[143],S[220],C[220]);
  fa FA_00000221 (C[177],S[143],C[144],S[221],C[221]);
  fa FA_00000222 (C[178],S[144],C[145],S[222],C[222]);
  fa FA_00000223 (C[179],S[145],C[146],S[223],C[223]);
  fa FA_00000224 (C[180],S[146],C[147],S[224],C[224]);
  fa FA_00000225 (C[181],S[147],C[148],S[225],C[225]);
  fa FA_00000226 (C[182],S[148],C[149],S[226],C[226]);
  fa FA_00000227 (C[183],S[149],C[150],S[227],C[227]);
  fa FA_00000228 (C[184],S[150],C[151],S[228],C[228]);
  fa FA_00000229 (C[185],S[151],C[152],S[229],C[229]);
  fa FA_00000230 (C[186],S[152],C[153],S[230],C[230]);
  fa FA_00000231 (C[187],S[153],C[154],S[231],C[231]);
  ha HA_00000232 (C[188],S[154],S[232],C[232]);
  ha HA_00000233 (C[189],C[84],S[233],C[233]);
  ha HA_00000234 (S[68],S[218],S[234],C[234]);
  ha HA_00000235 (S[174],S[219],S[235],C[235]);
  ha HA_00000236 (S[175],S[220],S[236],C[236]);
  ha HA_00000237 (S[176],S[221],S[237],C[237]);
  fa FA_00000238 (S[177],C[194],S[222],S[238],C[238]);
  fa FA_00000239 (S[194],C[195],S[223],S[239],C[239]);
  fa FA_00000240 (S[195],C[196],S[224],S[240],C[240]);
  fa FA_00000241 (S[196],C[197],S[225],S[241],C[241]);
  fa FA_00000242 (S[197],C[198],S[226],S[242],C[242]);
  fa FA_00000243 (S[198],C[199],S[227],S[243],C[243]);
  fa FA_00000244 (S[199],C[200],S[228],S[244],C[244]);
  fa FA_00000245 (S[200],C[201],S[229],S[245],C[245]);
  fa FA_00000246 (S[201],C[202],S[230],S[246],C[246]);
  fa FA_00000247 (S[202],C[203],S[231],S[247],C[247]);
  fa FA_00000248 (S[203],C[204],S[232],S[248],C[248]);
  fa FA_00000249 (S[204],C[205],S[233],S[249],C[249]);
  fa FA_00000250 (S[205],C[206],C[190],S[250],C[250]);
  fa FA_00000251 (S[206],C[207],C[191],S[251],C[251]);
  fa FA_00000252 (S[207],C[208],C[192],S[252],C[252]);
  fa FA_00000253 (S[208],C[209],C[193],S[253],C[253]);
  ha HA_00000254 (S[209],C[210],S[254],C[254]);
  ha HA_00000255 (S[210],C[211],S[255],C[255]);
  ha HA_00000256 (S[211],C[212],S[256],C[256]);
  ha HA_00000257 (S[212],C[213],S[257],C[257]);
  ha HA_00000258 (S[213],C[214],S[258],C[258]);
  ha HA_00000259 (S[215],C[216],S[259],C[259]);
  ha HA_00000260 (S[216],C[217],S[260],C[260]);
  fa FA_00000261 (S[217],C[234],C[218],S[261],C[261]);
  fa FA_00000262 (S[234],C[235],C[219],S[262],C[262]);
  fa FA_00000263 (S[235],C[236],C[220],S[263],C[263]);
  fa FA_00000264 (S[236],C[237],C[221],S[264],C[264]);
  fa FA_00000265 (S[237],C[238],C[222],S[265],C[265]);
  fa FA_00000266 (S[238],C[239],C[223],S[266],C[266]);
  fa FA_00000267 (S[239],C[240],C[224],S[267],C[267]);
  fa FA_00000268 (S[240],C[241],C[225],S[268],C[268]);
  fa FA_00000269 (S[241],C[242],C[226],S[269],C[269]);
  fa FA_00000270 (S[242],C[243],C[227],S[270],C[270]);
  fa FA_00000271 (S[243],C[244],C[228],S[271],C[271]);
  fa FA_00000272 (S[244],C[245],C[229],S[272],C[272]);
  fa FA_00000273 (S[245],C[246],C[230],S[273],C[273]);
  fa FA_00000274 (S[246],C[247],C[231],S[274],C[274]);
  fa FA_00000275 (S[247],C[248],C[232],S[275],C[275]);
  fa FA_00000276 (S[248],C[249],C[233],S[276],C[276]);
  ha HA_00000277 (S[249],C[250],S[277],C[277]);
  ha HA_00000278 (S[250],C[251],S[278],C[278]);
  ha HA_00000279 (S[251],C[252],S[279],C[279]);
  ha HA_00000280 (S[252],C[253],S[280],C[280]);
  ha HA_00000281 (S[253],C[254],S[281],C[281]);
  ha HA_00000282 (S[254],C[255],S[282],C[282]);
  ha HA_00000283 (S[255],C[256],S[283],C[283]);
  ha HA_00000284 (S[256],C[257],S[284],C[284]);
  ha HA_00000285 (S[257],C[258],S[285],C[285]);
  ha HA_00000286 (P[0][13],P[1][12],S[0],C[0]);
  fa FA_00000287 (P[0][14],P[1][13],P[2][12],S[1],C[1]);
  ha HA_00000288 (P[3][11],P[4][10],S[2],C[2]);
  fa FA_00000289 (P[0][15],P[1][14],P[2][13],S[3],C[3]);
  fa FA_00000290 (P[3][12],P[4][11],P[5][10],S[4],C[4]);
  ha HA_00000291 (P[6][9],P[7][8],S[5],C[5]);
  fa FA_00000292 (P[0][16],P[1][15],P[2][14],S[6],C[6]);
  fa FA_00000293 (P[3][13],P[4][12],P[5][11],S[7],C[7]);
  fa FA_00000294 (P[6][10],P[7][9],P[8][8],S[8],C[8]);
  ha HA_00000295 (P[9][7],P[10][6],S[9],C[9]);
  fa FA_00000296 (P[1][16],P[2][15],P[3][14],S[10],C[10]);
  fa FA_00000297 (P[4][13],P[5][12],P[6][11],S[11],C[11]);
  fa FA_00000298 (P[7][10],P[8][9],P[9][8],S[12],C[12]);
  ha HA_00000299 (P[10][7],P[11][6],S[13],C[13]);
  fa FA_00000300 (P[2][16],P[3][15],P[4][14],S[14],C[14]);
  fa FA_00000301 (P[5][13],P[6][12],P[7][11],S[15],C[15]);
  fa FA_00000302 (P[8][10],P[9][9],P[10][8],S[16],C[16]);
  fa FA_00000303 (P[3][16],P[4][15],P[5][14],S[17],C[17]);
  fa FA_00000304 (P[6][13],P[7][12],P[8][11],S[18],C[18]);
  fa FA_00000305 (P[4][16],P[5][15],P[6][14],S[19],C[19]);
  ha HA_00000306 (P[0][9],P[1][8],S[20],C[20]);
  fa FA_00000307 (P[0][10],P[1][9],P[2][8],S[21],C[21]);
  ha HA_00000308 (P[3][7],P[4][6],S[22],C[22]);
  fa FA_00000309 (P[0][11],P[1][10],P[2][9],S[23],C[23]);
  fa FA_00000310 (P[3][8],P[4][7],P[5][6],S[24],C[24]);
  ha HA_00000311 (P[6][5],P[7][4],S[25],C[25]);
  fa FA_00000312 (P[0][12],P[1][11],P[2][10],S[26],C[26]);
  fa FA_00000313 (P[3][9],P[4][8],P[5][7],S[27],C[27]);
  fa FA_00000314 (P[6][6],P[7][5],P[8][4],S[28],C[28]);
  ha HA_00000315 (P[9][3],P[10][2],S[29],C[29]);
  fa FA_00000316 (S[0],P[2][11],P[3][10],S[30],C[30]);
  fa FA_00000317 (P[4][9],P[5][8],P[6][7],S[31],C[31]);
  fa FA_00000318 (P[7][6],P[8][5],P[9][4],S[32],C[32]);
  fa FA_00000319 (P[10][3],P[11][2],P[12][1],S[33],C[33]);
  fa FA_00000320 (S[1],C[0],S[2],S[34],C[34]);
  fa FA_00000321 (P[5][9],P[6][8],P[7][7],S[35],C[35]);
  fa FA_00000322 (P[8][6],P[9][5],P[10][4],S[36],C[36]);
  fa FA_00000323 (P[11][3],P[12][2],P[13][1],S[37],C[37]);
  fa FA_00000324 (S[3],C[1],S[4],S[38],C[38]);
  fa FA_00000325 (C[2],S[5],P[8][7],S[39],C[39]);
  fa FA_00000326 (P[9][6],P[10][5],P[11][4],S[40],C[40]);
  fa FA_00000327 (P[12][3],P[13][2],P[14][1],S[41],C[41]);
  fa FA_00000328 (S[6],C[3],S[7],S[42],C[42]);
  fa FA_00000329 (C[4],S[8],C[5],S[43],C[43]);
  fa FA_00000330 (S[9],P[11][5],P[12][4],S[44],C[44]);
  fa FA_00000331 (P[13][3],P[14][2],P[15][1],S[45],C[45]);
  fa FA_00000332 (S[10],C[6],S[11],S[46],C[46]);
  fa FA_00000333 (C[7],S[12],C[8],S[47],C[47]);
  fa FA_00000334 (S[13],C[9],P[12][5],S[48],C[48]);
  fa FA_00000335 (P[13][4],P[14][3],P[15][2],S[49],C[49]);
  fa FA_00000336 (S[14],C[10],S[15],S[50],C[50]);
  fa FA_00000337 (C[11],S[16],C[12],S[51],C[51]);
  fa FA_00000338 (C[13],P[11][7],P[12][6],S[52],C[52]);
  fa FA_00000339 (P[13][5],P[14][4],P[15][3],S[53],C[53]);
  fa FA_00000340 (S[17],C[14],S[18],S[54],C[54]);
  fa FA_00000341 (C[15],C[16],P[9][10],S[55],C[55]);
  fa FA_00000342 (P[10][9],P[11][8],P[12][7],S[56],C[56]);
  fa FA_00000343 (P[13][6],P[14][5],P[15][4],S[57],C[57]);
  fa FA_00000344 (S[19],C[17],C[18],S[58],C[58]);
  fa FA_00000345 (P[7][13],P[8][12],P[9][11],S[59],C[59]);
  fa FA_00000346 (P[10][10],P[11][9],P[12][8],S[60],C[60]);
  fa FA_00000347 (P[13][7],P[14][6],P[15][5],S[61],C[61]);
  fa FA_00000348 (C[19],P[5][16],P[6][15],S[62],C[62]);
  fa FA_00000349 (P[7][14],P[8][13],P[9][12],S[63],C[63]);
  fa FA_00000350 (P[10][11],P[11][10],P[12][9],S[64],C[64]);
  fa FA_00000351 (P[13][8],P[14][7],P[15][6],S[65],C[65]);
  fa FA_00000352 (P[6][16],P[7][15],P[8][14],S[66],C[66]);
  fa FA_00000353 (P[9][13],P[10][12],P[11][11],S[67],C[67]);
  fa FA_00000354 (P[12][10],P[13][9],P[14][8],S[68],C[68]);
  fa FA_00000355 (P[7][16],P[8][15],P[9][14],S[69],C[69]);
  fa FA_00000356 (P[10][13],P[11][12],P[12][11],S[70],C[70]);
  fa FA_00000357 (P[8][16],P[9][15],P[10][14],S[71],C[71]);
  ha HA_00000358 (P[0][6],P[1][5],S[72],C[72]);
  fa FA_00000359 (P[0][7],P[1][6],P[2][5],S[73],C[73]);
  ha HA_00000360 (P[3][4],P[4][3],S[74],C[74]);
  fa FA_00000361 (P[0][8],P[1][7],P[2][6],S[75],C[75]);
  fa FA_00000362 (P[3][5],P[4][4],P[5][3],S[76],C[76]);
  ha HA_00000363 (P[6][2],P[7][1],S[77],C[77]);
  fa FA_00000364 (S[20],P[2][7],P[3][6],S[78],C[78]);
  fa FA_00000365 (P[4][5],P[5][4],P[6][3],S[79],C[79]);
  fa FA_00000366 (P[7][2],P[8][1],P[9][0],S[80],C[80]);
  fa FA_00000367 (S[21],C[20],S[22],S[81],C[81]);
  fa FA_00000368 (P[5][5],P[6][4],P[7][3],S[82],C[82]);
  fa FA_00000369 (P[8][2],P[9][1],P[10][0],S[83],C[83]);
  fa FA_00000370 (S[23],C[21],S[24],S[84],C[84]);
  fa FA_00000371 (C[22],S[25],P[8][3],S[85],C[85]);
  fa FA_00000372 (P[9][2],P[10][1],P[11][0],S[86],C[86]);
  fa FA_00000373 (S[26],C[23],S[27],S[87],C[87]);
  fa FA_00000374 (C[24],S[28],C[25],S[88],C[88]);
  fa FA_00000375 (S[29],P[11][1],P[12][0],S[89],C[89]);
  fa FA_00000376 (S[30],C[26],S[31],S[90],C[90]);
  fa FA_00000377 (C[27],S[32],C[28],S[91],C[91]);
  fa FA_00000378 (S[33],C[29],P[13][0],S[92],C[92]);
  fa FA_00000379 (S[34],C[30],S[35],S[93],C[93]);
  fa FA_00000380 (C[31],S[36],C[32],S[94],C[94]);
  fa FA_00000381 (S[37],C[33],P[14][0],S[95],C[95]);
  fa FA_00000382 (S[38],C[34],S[39],S[96],C[96]);
  fa FA_00000383 (C[35],S[40],C[36],S[97],C[97]);
  fa FA_00000384 (S[41],C[37],P[15][0],S[98],C[98]);
  fa FA_00000385 (S[42],C[38],S[43],S[99],C[99]);
  fa FA_00000386 (C[39],S[44],C[40],S[100],C[100]);
  fa FA_00000387 (S[45],C[41],P[16][0],S[101],C[101]);
  fa FA_00000388 (S[46],C[42],S[47],S[102],C[102]);
  fa FA_00000389 (C[43],S[48],C[44],S[103],C[103]);
  fa FA_00000390 (S[49],C[45],P[16][1],S[104],C[104]);
  fa FA_00000391 (S[50],C[46],S[51],S[105],C[105]);
  fa FA_00000392 (C[47],S[52],C[48],S[106],C[106]);
  fa FA_00000393 (S[53],C[49],P[16][2],S[107],C[107]);
  fa FA_00000394 (S[54],C[50],S[55],S[108],C[108]);
  fa FA_00000395 (C[51],S[56],C[52],S[109],C[109]);
  fa FA_00000396 (S[57],C[53],P[16][3],S[110],C[110]);
  fa FA_00000397 (S[58],C[54],S[59],S[111],C[111]);
  fa FA_00000398 (C[55],S[60],C[56],S[112],C[112]);
  fa FA_00000399 (S[61],C[57],P[16][4],S[113],C[113]);
  fa FA_00000400 (S[62],C[58],S[63],S[114],C[114]);
  fa FA_00000401 (C[59],S[64],C[60],S[115],C[115]);
  fa FA_00000402 (S[65],C[61],P[16][5],S[116],C[116]);
  fa FA_00000403 (S[66],C[62],S[67],S[117],C[117]);
  fa FA_00000404 (C[63],S[68],C[64],S[118],C[118]);
  fa FA_00000405 (C[65],P[15][7],P[16][6],S[119],C[119]);
  fa FA_00000406 (S[69],C[66],S[70],S[120],C[120]);
  fa FA_00000407 (C[67],C[68],P[13][10],S[121],C[121]);
  fa FA_00000408 (P[14][9],P[15][8],P[16][7],S[122],C[122]);
  fa FA_00000409 (S[71],C[69],C[70],S[123],C[123]);
  fa FA_00000410 (P[11][13],P[12][12],P[13][11],S[124],C[124]);
  fa FA_00000411 (P[14][10],P[15][9],P[16][8],S[125],C[125]);
  fa FA_00000412 (C[71],P[9][16],P[10][15],S[126],C[126]);
  fa FA_00000413 (P[11][14],P[12][13],P[13][12],S[127],C[127]);
  fa FA_00000414 (P[14][11],P[15][10],P[16][9],S[128],C[128]);
  fa FA_00000415 (P[10][16],P[11][15],P[12][14],S[129],C[129]);
  fa FA_00000416 (P[13][13],P[14][12],P[15][11],S[130],C[130]);
  fa FA_00000417 (P[11][16],P[12][15],P[13][14],S[131],C[131]);
  ha HA_00000418 (P[0][4],P[1][3],S[132],C[132]);
  fa FA_00000419 (P[0][5],P[1][4],P[2][3],S[133],C[133]);
  ha HA_00000420 (P[3][2],P[4][1],S[134],C[134]);
  fa FA_00000421 (S[72],P[2][4],P[3][3],S[135],C[135]);
  fa FA_00000422 (P[4][2],P[5][1],P[6][0],S[136],C[136]);
  fa FA_00000423 (S[73],C[72],S[74],S[137],C[137]);
  fa FA_00000424 (P[5][2],P[6][1],P[7][0],S[138],C[138]);
  fa FA_00000425 (S[75],C[73],S[76],S[139],C[139]);
  fa FA_00000426 (C[74],S[77],P[8][0],S[140],C[140]);
  fa FA_00000427 (S[78],C[75],S[79],S[141],C[141]);
  fa FA_00000428 (C[76],S[80],C[77],S[142],C[142]);
  fa FA_00000429 (S[81],C[78],S[82],S[143],C[143]);
  fa FA_00000430 (C[79],S[83],C[80],S[144],C[144]);
  fa FA_00000431 (S[84],C[81],S[85],S[145],C[145]);
  fa FA_00000432 (C[82],S[86],C[83],S[146],C[146]);
  fa FA_00000433 (S[87],C[84],S[88],S[147],C[147]);
  fa FA_00000434 (C[85],S[89],C[86],S[148],C[148]);
  fa FA_00000435 (S[90],C[87],S[91],S[149],C[149]);
  fa FA_00000436 (C[88],S[92],C[89],S[150],C[150]);
  fa FA_00000437 (S[93],C[90],S[94],S[151],C[151]);
  fa FA_00000438 (C[91],S[95],C[92],S[152],C[152]);
  fa FA_00000439 (S[96],C[93],S[97],S[153],C[153]);
  fa FA_00000440 (C[94],S[98],C[95],S[154],C[154]);
  fa FA_00000441 (S[99],C[96],S[100],S[155],C[155]);
  fa FA_00000442 (C[97],S[101],C[98],S[156],C[156]);
  fa FA_00000443 (S[102],C[99],S[103],S[157],C[157]);
  fa FA_00000444 (C[100],S[104],C[101],S[158],C[158]);
  fa FA_00000445 (S[105],C[102],S[106],S[159],C[159]);
  fa FA_00000446 (C[103],S[107],C[104],S[160],C[160]);
  fa FA_00000447 (S[108],C[105],S[109],S[161],C[161]);
  fa FA_00000448 (C[106],S[110],C[107],S[162],C[162]);
  fa FA_00000449 (S[111],C[108],S[112],S[163],C[163]);
  fa FA_00000450 (C[109],S[113],C[110],S[164],C[164]);
  fa FA_00000451 (S[114],C[111],S[115],S[165],C[165]);
  fa FA_00000452 (C[112],S[116],C[113],S[166],C[166]);
  fa FA_00000453 (S[117],C[114],S[118],S[167],C[167]);
  fa FA_00000454 (C[115],S[119],C[116],S[168],C[168]);
  fa FA_00000455 (S[120],C[117],S[121],S[169],C[169]);
  fa FA_00000456 (C[118],S[122],C[119],S[170],C[170]);
  fa FA_00000457 (S[123],C[120],S[124],S[171],C[171]);
  fa FA_00000458 (C[121],S[125],C[122],S[172],C[172]);
  fa FA_00000459 (S[126],C[123],S[127],S[173],C[173]);
  fa FA_00000460 (C[124],S[128],C[125],S[174],C[174]);
  fa FA_00000461 (S[129],C[126],S[130],S[175],C[175]);
  fa FA_00000462 (C[127],C[128],P[16][10],S[176],C[176]);
  fa FA_00000463 (S[131],C[129],C[130],S[177],C[177]);
  fa FA_00000464 (P[14][13],P[15][12],P[16][11],S[178],C[178]);
  fa FA_00000465 (C[131],P[12][16],P[13][15],S[179],C[179]);
  fa FA_00000466 (P[14][14],P[15][13],P[16][12],S[180],C[180]);
  fa FA_00000467 (P[13][16],P[14][15],P[15][14],S[181],C[181]);
  ha HA_00000468 (P[0][3],P[1][2],S[182],C[182]);
  fa FA_00000469 (S[132],P[2][2],P[3][1],S[183],C[183]);
  fa FA_00000470 (S[133],C[132],S[134],S[184],C[184]);
  fa FA_00000471 (S[135],C[133],S[136],S[185],C[185]);
  fa FA_00000472 (S[137],C[135],S[138],S[186],C[186]);
  fa FA_00000473 (S[139],C[137],S[140],S[187],C[187]);
  fa FA_00000474 (S[141],C[139],S[142],S[188],C[188]);
  fa FA_00000475 (S[143],C[141],S[144],S[189],C[189]);
  fa FA_00000476 (S[145],C[143],S[146],S[190],C[190]);
  fa FA_00000477 (S[147],C[145],S[148],S[191],C[191]);
  fa FA_00000478 (S[149],C[147],S[150],S[192],C[192]);
  fa FA_00000479 (S[151],C[149],S[152],S[193],C[193]);
  fa FA_00000480 (S[153],C[151],S[154],S[194],C[194]);
  fa FA_00000481 (S[155],C[153],S[156],S[195],C[195]);
  fa FA_00000482 (S[157],C[155],S[158],S[196],C[196]);
  fa FA_00000483 (S[159],C[157],S[160],S[197],C[197]);
  fa FA_00000484 (S[161],C[159],S[162],S[198],C[198]);
  fa FA_00000485 (S[163],C[161],S[164],S[199],C[199]);
  fa FA_00000486 (S[165],C[163],S[166],S[200],C[200]);
  fa FA_00000487 (S[167],C[165],S[168],S[201],C[201]);
  fa FA_00000488 (S[169],C[167],S[170],S[202],C[202]);
  fa FA_00000489 (S[171],C[169],S[172],S[203],C[203]);
  fa FA_00000490 (S[173],C[171],S[174],S[204],C[204]);
  fa FA_00000491 (S[175],C[173],S[176],S[205],C[205]);
  fa FA_00000492 (S[177],C[175],S[178],S[206],C[206]);
  fa FA_00000493 (S[179],C[177],S[180],S[207],C[207]);
  fa FA_00000494 (S[181],C[179],C[180],S[208],C[208]);
  fa FA_00000495 (C[181],P[14][16],P[15][15],S[209],C[209]);
  ha HA_00000496 (P[0][2],P[1][1],S[210],C[210]);
  fa FA_00000497 (S[182],P[2][1],P[3][0],S[211],C[211]);
  fa FA_00000498 (S[183],C[182],P[4][0],S[212],C[212]);
  fa FA_00000499 (S[184],C[183],P[5][0],S[213],C[213]);
  fa FA_00000500 (S[185],C[184],C[134],S[214],C[214]);
  fa FA_00000501 (S[186],C[185],C[136],S[215],C[215]);
  fa FA_00000502 (S[187],C[186],C[138],S[216],C[216]);
  fa FA_00000503 (S[188],C[187],C[140],S[217],C[217]);
  fa FA_00000504 (S[189],C[188],C[142],S[218],C[218]);
  fa FA_00000505 (S[190],C[189],C[144],S[219],C[219]);
  fa FA_00000506 (S[191],C[190],C[146],S[220],C[220]);
  fa FA_00000507 (S[192],C[191],C[148],S[221],C[221]);
  fa FA_00000508 (S[193],C[192],C[150],S[222],C[222]);
  fa FA_00000509 (S[194],C[193],C[152],S[223],C[223]);
  fa FA_00000510 (S[195],C[194],C[154],S[224],C[224]);
  fa FA_00000511 (S[196],C[195],C[156],S[225],C[225]);
  fa FA_00000512 (S[197],C[196],C[158],S[226],C[226]);
  fa FA_00000513 (S[198],C[197],C[160],S[227],C[227]);
  fa FA_00000514 (S[199],C[198],C[162],S[228],C[228]);
  fa FA_00000515 (S[200],C[199],C[164],S[229],C[229]);
  fa FA_00000516 (S[201],C[200],C[166],S[230],C[230]);
  fa FA_00000517 (S[202],C[201],C[168],S[231],C[231]);
  fa FA_00000518 (S[203],C[202],C[170],S[232],C[232]);
  fa FA_00000519 (S[204],C[203],C[172],S[233],C[233]);
  fa FA_00000520 (S[205],C[204],C[174],S[234],C[234]);
  fa FA_00000521 (S[206],C[205],C[176],S[235],C[235]);
  fa FA_00000522 (S[207],C[206],C[178],S[236],C[236]);
  fa FA_00000523 (S[208],C[207],P[16][13],S[237],C[237]);
  fa FA_00000524 (S[209],C[208],P[16][14],S[238],C[238]);
  fa FA_00000525 (C[209],P[15][16],P[16][15],S[239],C[239]);

  assign z0[0] = P[0][0];
  assign z0[1] = P[0][1];
  assign z0[2] = S[210];
  assign z0[3] = S[211];
  assign z0[4] = S[212];
  assign z0[5] = S[213];
  assign z0[6] = S[214];
  assign z0[7] = S[215];
  assign z0[8] = S[216];
  assign z0[9] = S[217];
  assign z0[10] = S[218];
  assign z0[11] = S[219];
  assign z0[12] = S[220];
  assign z0[13] = S[221];
  assign z0[14] = S[222];
  assign z0[15] = S[223];
  assign z0[16] = S[224];
  assign z0[17] = S[225];
  assign z0[18] = S[226];
  assign z0[19] = S[227];
  assign z0[20] = S[228];
  assign z0[21] = S[229];
  assign z0[22] = S[230];
  assign z0[23] = S[231];
  assign z0[24] = S[232];
  assign z0[25] = S[233];
  assign z0[26] = S[234];
  assign z0[27] = S[235];
  assign z0[28] = S[236];
  assign z0[29] = S[237];
  assign z0[30] = S[238];
  assign z0[31] = S[239];
  assign z0[32] = C[239];
  assign z0[33] = 0;
  assign z1[0] = 0;
  assign z1[1] = P[1][0];
  assign z1[2] = P[2][0];
  assign z1[3] = C[210];
  assign z1[4] = C[211];
  assign z1[5] = C[212];
  assign z1[6] = C[213];
  assign z1[7] = C[214];
  assign z1[8] = C[215];
  assign z1[9] = C[216];
  assign z1[10] = C[217];
  assign z1[11] = C[218];
  assign z1[12] = C[219];
  assign z1[13] = C[220];
  assign z1[14] = C[221];
  assign z1[15] = C[222];
  assign z1[16] = C[223];
  assign z1[17] = C[224];
  assign z1[18] = C[225];
  assign z1[19] = C[226];
  assign z1[20] = C[227];
  assign z1[21] = C[228];
  assign z1[22] = C[229];
  assign z1[23] = C[230];
  assign z1[24] = C[231];
  assign z1[25] = C[232];
  assign z1[26] = C[233];
  assign z1[27] = C[234];
  assign z1[28] = C[235];
  assign z1[29] = C[236];
  assign z1[30] = C[237];
  assign z1[31] = C[238];
  assign z1[32] = P[16][16];
  assign z1[33] = 0;

endmodule
